magic
tech sky130A
magscale 1 2
timestamp 1671181216
<< obsli1 >>
rect 1104 2159 28888 31569
<< obsm1 >>
rect 566 2128 29048 31600
<< metal2 >>
rect 570 33200 626 34000
rect 1674 33200 1730 34000
rect 2778 33200 2834 34000
rect 3882 33200 3938 34000
rect 4986 33200 5042 34000
rect 6090 33200 6146 34000
rect 7194 33200 7250 34000
rect 8298 33200 8354 34000
rect 9402 33200 9458 34000
rect 10506 33200 10562 34000
rect 11610 33200 11666 34000
rect 12714 33200 12770 34000
rect 13818 33200 13874 34000
rect 14922 33200 14978 34000
rect 16026 33200 16082 34000
rect 17130 33200 17186 34000
rect 18234 33200 18290 34000
rect 19338 33200 19394 34000
rect 20442 33200 20498 34000
rect 21546 33200 21602 34000
rect 22650 33200 22706 34000
rect 23754 33200 23810 34000
rect 24858 33200 24914 34000
rect 25962 33200 26018 34000
rect 27066 33200 27122 34000
rect 28170 33200 28226 34000
rect 29274 33200 29330 34000
<< obsm2 >>
rect 682 33144 1618 33200
rect 1786 33144 2722 33200
rect 2890 33144 3826 33200
rect 3994 33144 4930 33200
rect 5098 33144 6034 33200
rect 6202 33144 7138 33200
rect 7306 33144 8242 33200
rect 8410 33144 9346 33200
rect 9514 33144 10450 33200
rect 10618 33144 11554 33200
rect 11722 33144 12658 33200
rect 12826 33144 13762 33200
rect 13930 33144 14866 33200
rect 15034 33144 15970 33200
rect 16138 33144 17074 33200
rect 17242 33144 18178 33200
rect 18346 33144 19282 33200
rect 19450 33144 20386 33200
rect 20554 33144 21490 33200
rect 21658 33144 22594 33200
rect 22762 33144 23698 33200
rect 23866 33144 24802 33200
rect 24970 33144 25906 33200
rect 26074 33144 27010 33200
rect 27178 33144 28114 33200
rect 28282 33144 29042 33200
rect 572 2139 29042 33144
<< metal3 >>
rect 29200 31832 30000 31952
rect 29200 31152 30000 31272
rect 0 30880 800 31000
rect 29200 30472 30000 30592
rect 0 30200 800 30320
rect 29200 29792 30000 29912
rect 0 29520 800 29640
rect 29200 29112 30000 29232
rect 0 28840 800 28960
rect 29200 28432 30000 28552
rect 0 28160 800 28280
rect 29200 27752 30000 27872
rect 0 27480 800 27600
rect 29200 27072 30000 27192
rect 0 26800 800 26920
rect 29200 26392 30000 26512
rect 0 26120 800 26240
rect 29200 25712 30000 25832
rect 0 25440 800 25560
rect 29200 25032 30000 25152
rect 0 24760 800 24880
rect 29200 24352 30000 24472
rect 0 24080 800 24200
rect 29200 23672 30000 23792
rect 0 23400 800 23520
rect 29200 22992 30000 23112
rect 0 22720 800 22840
rect 29200 22312 30000 22432
rect 0 22040 800 22160
rect 29200 21632 30000 21752
rect 0 21360 800 21480
rect 29200 20952 30000 21072
rect 0 20680 800 20800
rect 29200 20272 30000 20392
rect 0 20000 800 20120
rect 29200 19592 30000 19712
rect 0 19320 800 19440
rect 29200 18912 30000 19032
rect 0 18640 800 18760
rect 29200 18232 30000 18352
rect 0 17960 800 18080
rect 29200 17552 30000 17672
rect 0 17280 800 17400
rect 29200 16872 30000 16992
rect 0 16600 800 16720
rect 29200 16192 30000 16312
rect 0 15920 800 16040
rect 29200 15512 30000 15632
rect 0 15240 800 15360
rect 29200 14832 30000 14952
rect 0 14560 800 14680
rect 29200 14152 30000 14272
rect 0 13880 800 14000
rect 29200 13472 30000 13592
rect 0 13200 800 13320
rect 29200 12792 30000 12912
rect 0 12520 800 12640
rect 29200 12112 30000 12232
rect 0 11840 800 11960
rect 29200 11432 30000 11552
rect 0 11160 800 11280
rect 29200 10752 30000 10872
rect 0 10480 800 10600
rect 29200 10072 30000 10192
rect 0 9800 800 9920
rect 29200 9392 30000 9512
rect 0 9120 800 9240
rect 29200 8712 30000 8832
rect 0 8440 800 8560
rect 29200 8032 30000 8152
rect 0 7760 800 7880
rect 29200 7352 30000 7472
rect 0 7080 800 7200
rect 29200 6672 30000 6792
rect 0 6400 800 6520
rect 29200 5992 30000 6112
rect 0 5720 800 5840
rect 29200 5312 30000 5432
rect 0 5040 800 5160
rect 29200 4632 30000 4752
rect 0 4360 800 4480
rect 29200 3952 30000 4072
rect 0 3680 800 3800
rect 29200 3272 30000 3392
rect 0 3000 800 3120
rect 29200 2592 30000 2712
rect 29200 1912 30000 2032
<< obsm3 >>
rect 800 31752 29120 31925
rect 800 31352 29378 31752
rect 800 31080 29120 31352
rect 880 31072 29120 31080
rect 880 30800 29378 31072
rect 800 30672 29378 30800
rect 800 30400 29120 30672
rect 880 30392 29120 30400
rect 880 30120 29378 30392
rect 800 29992 29378 30120
rect 800 29720 29120 29992
rect 880 29712 29120 29720
rect 880 29440 29378 29712
rect 800 29312 29378 29440
rect 800 29040 29120 29312
rect 880 29032 29120 29040
rect 880 28760 29378 29032
rect 800 28632 29378 28760
rect 800 28360 29120 28632
rect 880 28352 29120 28360
rect 880 28080 29378 28352
rect 800 27952 29378 28080
rect 800 27680 29120 27952
rect 880 27672 29120 27680
rect 880 27400 29378 27672
rect 800 27272 29378 27400
rect 800 27000 29120 27272
rect 880 26992 29120 27000
rect 880 26720 29378 26992
rect 800 26592 29378 26720
rect 800 26320 29120 26592
rect 880 26312 29120 26320
rect 880 26040 29378 26312
rect 800 25912 29378 26040
rect 800 25640 29120 25912
rect 880 25632 29120 25640
rect 880 25360 29378 25632
rect 800 25232 29378 25360
rect 800 24960 29120 25232
rect 880 24952 29120 24960
rect 880 24680 29378 24952
rect 800 24552 29378 24680
rect 800 24280 29120 24552
rect 880 24272 29120 24280
rect 880 24000 29378 24272
rect 800 23872 29378 24000
rect 800 23600 29120 23872
rect 880 23592 29120 23600
rect 880 23320 29378 23592
rect 800 23192 29378 23320
rect 800 22920 29120 23192
rect 880 22912 29120 22920
rect 880 22640 29378 22912
rect 800 22512 29378 22640
rect 800 22240 29120 22512
rect 880 22232 29120 22240
rect 880 21960 29378 22232
rect 800 21832 29378 21960
rect 800 21560 29120 21832
rect 880 21552 29120 21560
rect 880 21280 29378 21552
rect 800 21152 29378 21280
rect 800 20880 29120 21152
rect 880 20872 29120 20880
rect 880 20600 29378 20872
rect 800 20472 29378 20600
rect 800 20200 29120 20472
rect 880 20192 29120 20200
rect 880 19920 29378 20192
rect 800 19792 29378 19920
rect 800 19520 29120 19792
rect 880 19512 29120 19520
rect 880 19240 29378 19512
rect 800 19112 29378 19240
rect 800 18840 29120 19112
rect 880 18832 29120 18840
rect 880 18560 29378 18832
rect 800 18432 29378 18560
rect 800 18160 29120 18432
rect 880 18152 29120 18160
rect 880 17880 29378 18152
rect 800 17752 29378 17880
rect 800 17480 29120 17752
rect 880 17472 29120 17480
rect 880 17200 29378 17472
rect 800 17072 29378 17200
rect 800 16800 29120 17072
rect 880 16792 29120 16800
rect 880 16520 29378 16792
rect 800 16392 29378 16520
rect 800 16120 29120 16392
rect 880 16112 29120 16120
rect 880 15840 29378 16112
rect 800 15712 29378 15840
rect 800 15440 29120 15712
rect 880 15432 29120 15440
rect 880 15160 29378 15432
rect 800 15032 29378 15160
rect 800 14760 29120 15032
rect 880 14752 29120 14760
rect 880 14480 29378 14752
rect 800 14352 29378 14480
rect 800 14080 29120 14352
rect 880 14072 29120 14080
rect 880 13800 29378 14072
rect 800 13672 29378 13800
rect 800 13400 29120 13672
rect 880 13392 29120 13400
rect 880 13120 29378 13392
rect 800 12992 29378 13120
rect 800 12720 29120 12992
rect 880 12712 29120 12720
rect 880 12440 29378 12712
rect 800 12312 29378 12440
rect 800 12040 29120 12312
rect 880 12032 29120 12040
rect 880 11760 29378 12032
rect 800 11632 29378 11760
rect 800 11360 29120 11632
rect 880 11352 29120 11360
rect 880 11080 29378 11352
rect 800 10952 29378 11080
rect 800 10680 29120 10952
rect 880 10672 29120 10680
rect 880 10400 29378 10672
rect 800 10272 29378 10400
rect 800 10000 29120 10272
rect 880 9992 29120 10000
rect 880 9720 29378 9992
rect 800 9592 29378 9720
rect 800 9320 29120 9592
rect 880 9312 29120 9320
rect 880 9040 29378 9312
rect 800 8912 29378 9040
rect 800 8640 29120 8912
rect 880 8632 29120 8640
rect 880 8360 29378 8632
rect 800 8232 29378 8360
rect 800 7960 29120 8232
rect 880 7952 29120 7960
rect 880 7680 29378 7952
rect 800 7552 29378 7680
rect 800 7280 29120 7552
rect 880 7272 29120 7280
rect 880 7000 29378 7272
rect 800 6872 29378 7000
rect 800 6600 29120 6872
rect 880 6592 29120 6600
rect 880 6320 29378 6592
rect 800 6192 29378 6320
rect 800 5920 29120 6192
rect 880 5912 29120 5920
rect 880 5640 29378 5912
rect 800 5512 29378 5640
rect 800 5240 29120 5512
rect 880 5232 29120 5240
rect 880 4960 29378 5232
rect 800 4832 29378 4960
rect 800 4560 29120 4832
rect 880 4552 29120 4560
rect 880 4280 29378 4552
rect 800 4152 29378 4280
rect 800 3880 29120 4152
rect 880 3872 29120 3880
rect 880 3600 29378 3872
rect 800 3472 29378 3600
rect 800 3200 29120 3472
rect 880 3192 29120 3200
rect 880 2920 29378 3192
rect 800 2792 29378 2920
rect 800 2512 29120 2792
rect 800 2143 29378 2512
<< metal4 >>
rect 4417 2128 4737 31600
rect 7890 2128 8210 31600
rect 11363 2128 11683 31600
rect 14836 2128 15156 31600
rect 18309 2128 18629 31600
rect 21782 2128 22102 31600
rect 25255 2128 25575 31600
rect 28728 2128 29048 31600
<< labels >>
rlabel metal3 s 29200 1912 30000 2032 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 29200 22312 30000 22432 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 29200 24352 30000 24472 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 29200 26392 30000 26512 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 29200 28432 30000 28552 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 29200 30472 30000 30592 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 29274 33200 29330 34000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 25962 33200 26018 34000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 22650 33200 22706 34000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 19338 33200 19394 34000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 16026 33200 16082 34000 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 29200 3952 30000 4072 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 12714 33200 12770 34000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 9402 33200 9458 34000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 6090 33200 6146 34000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 2778 33200 2834 34000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 30880 800 31000 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 26800 800 26920 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 24760 800 24880 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 29200 5992 30000 6112 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 18640 800 18760 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 29200 8032 30000 8152 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 29200 10072 30000 10192 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 29200 12112 30000 12232 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 29200 14152 30000 14272 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 29200 16192 30000 16312 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 29200 18232 30000 18352 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 29200 20272 30000 20392 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 29200 3272 30000 3392 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 29200 23672 30000 23792 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 29200 25712 30000 25832 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 29200 27752 30000 27872 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 29200 29792 30000 29912 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 29200 31832 30000 31952 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 27066 33200 27122 34000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 23754 33200 23810 34000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 20442 33200 20498 34000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 17130 33200 17186 34000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 13818 33200 13874 34000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 29200 5312 30000 5432 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 10506 33200 10562 34000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 7194 33200 7250 34000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 3882 33200 3938 34000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 570 33200 626 34000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 29520 800 29640 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 27480 800 27600 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 25440 800 25560 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 23400 800 23520 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 29200 7352 30000 7472 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 17280 800 17400 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 13200 800 13320 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 9120 800 9240 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 29200 9392 30000 9512 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 29200 11432 30000 11552 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 29200 13472 30000 13592 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 29200 15512 30000 15632 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 29200 17552 30000 17672 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 29200 19592 30000 19712 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 29200 21632 30000 21752 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 29200 2592 30000 2712 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 29200 22992 30000 23112 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 29200 25032 30000 25152 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 29200 27072 30000 27192 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 29200 29112 30000 29232 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 29200 31152 30000 31272 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 28170 33200 28226 34000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 24858 33200 24914 34000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 21546 33200 21602 34000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 18234 33200 18290 34000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 14922 33200 14978 34000 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 29200 4632 30000 4752 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 11610 33200 11666 34000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 8298 33200 8354 34000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 4986 33200 5042 34000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 1674 33200 1730 34000 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 30200 800 30320 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 28160 800 28280 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 24080 800 24200 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 29200 6672 30000 6792 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 15920 800 16040 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 13880 800 14000 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 11840 800 11960 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 9800 800 9920 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 7760 800 7880 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 5720 800 5840 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 3680 800 3800 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 29200 8712 30000 8832 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 29200 10752 30000 10872 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 29200 12792 30000 12912 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 29200 14832 30000 14952 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 29200 16872 30000 16992 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 29200 18912 30000 19032 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 29200 20952 30000 21072 6 io_out[9]
port 114 nsew signal output
rlabel metal4 s 4417 2128 4737 31600 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 11363 2128 11683 31600 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 18309 2128 18629 31600 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 25255 2128 25575 31600 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 7890 2128 8210 31600 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 14836 2128 15156 31600 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 21782 2128 22102 31600 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 28728 2128 29048 31600 6 vssd1
port 116 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 34000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 502686
string GDS_FILE /home/runner/work/xls_workshop_tapeout_test_all_branch/xls_workshop_tapeout_test_all_branch/openlane/tiny_user_project/runs/22_12_16_08_58/results/signoff/tiny_user_project.magic.gds
string GDS_START 23768
<< end >>

